module ALU#(
    parameter WIDTH = 32,
    parameter REGBITS = 5,
)(
    input [5:0] opcode,
    input 
);







endmodule